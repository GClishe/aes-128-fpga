
// as of right now, I have no idea how the FPGA memory works. I do not yet know how I should setup the ports for this module
module vector_rom (

);